b0VIM 7.4      ���U�?l �  gangadhar                               Dev                                     ~gangadhar/erpnext/verve_wale/frappe-bench/apps/church_ministry/church_ministry/church_ministry/doctype/member/member.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           n                            l       o                     c       �                     \       >                    K       �                    L       �                    Z       1                    ^       �                    H       �                    -       0                           ]                    &       y             	       N       �             
       K       �                    M       8                    )       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     n       �  �  �  X  J  >    �  �  �  �  �  m  l  j  T  K  �  �  �  m  U  9  %  �  �  �  �  ^  E  (    �  �  �  �  _  D         �
  �
  �
  �
  q
  L
  =
  
  �	  �	  �	  �	  �	  �	  c	  >	  	  �  �  �  �  h  R  2  1  �  �  �  [  L  D  �  �  �  �  �  �  �  x  V    �  �  �  |  Y    �  �  �  z  ^  ]  \  <    �  (  %    �  t  s  `  4  �  �  �  �  �        ### web sevices   				frappe.throw(_('{0} is not a valid email id').format(doc.email_id)) 			if not validate_email_add(doc.email_id): 		if doc.email_id:  		# 		frappe.throw(_("When and Where is Mandatory if 'Baptisum Status' is 'Yes'..!")) 		# 	if not doc.baptism_when or not doc.baptism_where : 		# if doc.baptisum_status=='Yes': 		 			frappe.throw(_("Date of Joining '{0}' must be greater than Date of Birth '{1}'").format(doc.date_of_join, doc.date_of_birth)) 		if doc.date_of_birth and doc.date_of_join and getdate(doc.date_of_birth) >= getdate(doc.date_of_join):		 		#frappe.errprint("in date of birth ") def validate_birth(doc,method):   	return ' or '.join(cond)   		cond.append('region="%s"'%(filters.get('region'))) 	elif filters.get('region'): 		cond.append('zone="%s"'%(filters.get('zone'))) 	elif filters.get('zone'): 		cond.append('church_group="%s"'%(filters.get('church_group'))) 	elif filters.get('church_group'): 		cond.append('church="%s"'%(filters.get('church'))) 	elif filters.get('church'): 		cond.append('pcf="%s"'%(filters.get('pcf'))) 	elif filters.get('pcf'): 		cond.append('senior_cell="%s"'%(filters.get('senior_cell'))) 	elif filters.get('senior_cell'): 		cond.append('cell="%s"'%(filters.get('cell'))) 	if filters.get('cell'): 	cond=[] def get_conditions(filters):   		return value 		value=frappe.db.sql("select name from `tab%s`"%(filters.get('doctype'))) 	else : 		return value 		value=frappe.db.sql("select name from `tab%s` where %s"%(filters.get('doctype'),conditions)) 	if conditions: 	conditions=get_conditions(filters) def get_list(doctype, txt, searchfield, start, page_len, filters):  			self.user_id = self.email_id 			frappe.db.commit() 			frappe.db.sql("update `tabMember` set flag='SetPerm' where name='%s'"%(self.name)) 			v.insert() 			v.defvalue = self.name  			v.defkey = 'Member' 			v.parent = self.email_id 			v.parenttype = 'User Permission' 			v.parentfield = 'system_defaults' 			v = frappe.new_doc("DefaultValue") 			r.insert() 			r.role='Member' 			r.parenttype='User' 			r.parentfield='user_roles' 			r.parent=self.email_id 			r=frappe.new_doc("UserRole") 				frappe.flags.mute_emails = True 				u.insert() 				frappe.flags.mute_emails = False 				u.new_password = 'password' 				u.first_name = self.member_name 				u.email=self.email_id 				u = frappe.new_doc("User") 			if not usr_id:  			# 	perm = 'Churches' 			# 	r_user = 'Bible Study Class Teacher' 			# 	c_user = self.church 			# elif self.member_designation=='Bible Study Class Teacher': 			# 	perm = 'Member' 			# 	r_user = 'Member' 			# 	c_user = self.name 			# elif self.member_designation=='Member': 			# 	perm = 'Cells' 			# 	r_user = 'Cell Leader' 			# 	c_user = self.cell 			# elif self.member_designation=='Cell Leader': 			# 	perm = 'Senior Cells' 			# 	r_user = 'Senior Cell Leader' 			# 	c_user = self.senior_cell 			# elif self.member_designation=='Sr.Cell Leader': 			# 	perm = 'PCFs' 			# 	r_user = 'PCF Leader' 			# 	c_user = self.pcf 			# if  self.member_designation=='PCF Leader': 			# frappe.errprint("user creation") 		if self.flag=='not' and self.email_id: 		usr_id=frappe.db.sql("select name from `tabUser` where name='%s'"%(self.email_id),as_list=1) 		# pass 	def on_update(self): 	  class Member(Document):  from gcm import GCM  import base64 from frappe.utils import getdate, validate_email_add, cint,cstr,now from frappe import throw, _, msgprint from frappe.model.document import Document import json import frappe from __future__ import unicode_literals  # For license information, please see license.txt # Copyright (c) 2013, New Indictrans Technologies Pvt. Ltd. and contributors ad  �  �     )       �  �  �  �  �  �  �  `  X  1  )      �  P  3  !    �  �  �  �  G  �  �  V  @      �
  �
  �
  3
  *
  �	  �	  o	  X	  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            return "Successfully message has been sent"         frappe.sendmail(recipients=dts['recipents'], sender='verve@lws.com', content=dts['message'], subject='Message Broadcast') 	print "sending email"     if dts['email']: 		print "sending push notification"         	res = gcm.json_request(registration_ids=res, data=data,collapse_key='uptoyou', delay_while_idle=True, time_to_live=3600) 	if res: 	res=frappe.db.sql("select device_id from tabUser where name in ('%s')" % "','".join(map(str,rc_list)),as_list=1) 	gcm = GCM('AIzaSyBIc4LYCnUU9wFV_pBoFHHzLoGm_xHl-5k') 	data['Message']=dts['message'] 	data={}     if dts['push']:     rc_list=dts['recipents'].split(',') 		print "sending sms"     		send_sms([ x[0] for x in rc_list ], cstr(dts['message']))     	if rc_list: 	rc_list=frappe.db.sql("select phone_1 from tabMember where phone_1 is not null and email_id in ('%s')" %(dts['recipents'].replace(",","','")),as_list=1)               from erpnext.setup.doctype.sms_settings.sms_settings import send_sms     if dts['sms']:         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     from frappe.model.db_query import DatabaseQuery     #print dts     dts=json.loads(data)     """     this will return recipents details     """ def message_braudcast_send(data): @frappe.whitelist(allow_guest=True)       return res     #print res     res=frappe.db.sql(qry,as_dict=1)         qry="select name,member_name as ftv_name,email_id,phone_1 from tabMember where email_id in (select distinct parent from tabUserRole where role in ('PCF Leader','Cell Leader','Senior Cell Leader','Church Pastor','Group Church Pastor','Regional Pastor','Zonal Pastor'))" ad  �   5     ^       �  j  M  ;  *  
  �  �  �  w  W  �  �  �  �  �  �  o  V  �  �  �  �  �  k  ,  "    �  �  `  1  	  �
  �
  �
  U
  F
  E
  D
   
  
  �	  �	  f	  I	  7	  &	  	  �  �  �  �  l  K      �  �  �  �  �  o  P  (    �  �  �  �  �  k  B    �  �  �  ^  O  N  M  L  (    �  }  `  N  =    �  �  F  5                                                                                                                                                                           #print(data)     #data=frappe.db.sql("""select name ,owner as assignee,subject ,exp_end_date,status,priority,description,replace(replace(replace(SUBSTRING_INDEX(_assign,',',1),'"',''),'[',''),']','') as _assign,cell,senior_cell,pcf from `tabTask` where status in ('Open','Working' ) and exp_start_date is not null and owner='%s' or _assign like '%%%s%%' """ %(dts['username'],dts['username']),as_dict=True)         }                     "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def task_list(data): @frappe.whitelist(allow_guest=True)        return res     res=frappe.db.sql("select name from `tab%s` where %s='%s'"  %(fields[fieldname],wheres[tablename],dts['name']),as_dict=True)     fieldname=dts['tbl']     }             "Regions":"Zones"             "Zones":"Group Churches",             "Group Churches":"Churches",             "Churches":"PCFs",             "PCFs":"Senior Cells",             "Senior Cells":"Cells",     fields={     #}     #        "Regions":"zone"     #        "Zones":"church_group",     #        "Group Churches":"church",     #        "Churches":"pcf",     #        "PCFs":"senior_cell",     #        "Senior Cells":"name",     #fields={     tablename=dts['tbl']     }             "Regions":"region"             "Zones":"zone",             "Group Churches":"church_group",             "Churches":"church",             "PCFs":"pcf",             "Senior Cells":"senior_cell",     wheres={         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     #print dts     dts=json.loads(data) def get_lists(data): @frappe.whitelist(allow_guest=True)       return res     res=frappe.db.sql("select %s from `tab%s` where name='%s'"  %(dictnory[tablename],dts['tbl'],dts['name']),as_dict=True)     tablename=dts['tbl']     }         "Zones":"region"         "Group Churches":"zone,region",         "Churches":"church_group,zone,region",         "PCFs":"church,church_group,zone,region",         "Senior Cells":"pcf,church,church_group,zone,region",         "Cells":"senior_cell,pcf,church,church_group,zone,region",     dictnory={         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     print dts     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def get_hierarchy(data): @frappe.whitelist(allow_guest=True)        return "Updated Your Event Attendance"         frappe.db.sql("update `tabEvent Attendace Details` set present=%s where name=%s",(record['present'],record['name']))             record['present']=0         if not record['present'] :     for record in dts['records']:         }                      "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) ad     R     H       z  j  i  h  D  *    �  w  e  T  4  �  �  �  �  
  �	  �	  �	  �	  �	  *	  	  �  �  �  �  }  j  M  )    �  �  �  �  W  �  A  7  �  Y  X  4      �  i  W  F  &  �  �  S  C  B  A      �  p  S  A  0    �  �  �  �  j  R  Q                            del dts['assignee']     dts['owner']=dts['username']     dts['doctype']='Task'     dts['exp_start_date']=now()         }                   "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def create_task(data): @frappe.whitelist(allow_guest=True)       return data     data=frappe.db.sql("select a.member_name from tabMember a,tabUser b where a.user_id=b.name and a.cell=%s",dts['cell'],as_dict=True)         }                   "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def cell_members(data): @frappe.whitelist(allow_guest=True)          return "Task Details updated Successfully"         frappe.db.sql("update `tabTask` set description=%s,status=%s,_assign=%s where name=%s",(dts['description'],dts['status'],dts['_assign'],dts['name']),as_dict=True)     else:         return "Created followup taks "+ma.name+" and closed old task "+dts['name']         frappe.db.sql("update `tabTask` set description=%s,status='Closed',closing_date=%s where name=%s",('Closed the task and created followup task '+ma.name ,now(),dts['name']),as_dict=True)         ma.insert(ignore_permissions=True)         ma = frappe.get_doc(dts) 	del dts['_assign']         del dts['assignee']         dts['subject']='followup task for '+dts['name']         dts['doctype']='Task'         dts['exp_start_date']=now()     if dts['followup_task']:         }                          "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     print dts     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def task_update(data): @frappe.whitelist(allow_guest=True)      return data     data=frappe.db.sql("""select  a.name ,b.owner as _assign,b.assigned_by as assignee,a.subject ,a.exp_end_date,a.status,a.priority,a.description,a.cell,a.senior_cell,a.pcf from `tabTask` a, `tabToDo` b where a.status in ('Open','Working' )  and a.name=b.reference_name and a.exp_start_date is not null and a.owner='%s' or b.assigned_by='%s' """ %(dts['username'],dts['username']),as_dict=True)     #rint(data)     #ata=frappe.db.sql("""select name ,owner as assignee,subject ,exp_end_date,status,priority,description,replace(replace(replace(SUBSTRING_INDEX(_assign,',',1),'"',''),'[',''),']','') as _assign,cell,senior_cell,pcf from `tabTask` where status in ('Open','Working' ) and exp_start_date is not null """ ,as_dict=True)         }                     "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def task_list_team(data): @frappe.whitelist(allow_guest=True)       return data     data=frappe.db.sql("""select  a.name ,b.owner as _assign,b.assigned_by as assignee,a.subject ,a.exp_end_date,a.status,a.priority,a.description,a.cell,a.senior_cell,a.pcf from `tabTask` a, `tabToDo` b where a.status in ('Open','Working' )  and a.name=b.reference_name and a.exp_start_date is not null and a.owner='%s' or _assign='%s' """ %(dts['username'],dts['username']),as_dict=True) ad  :   
     -       �  �  �  }  |  {  z  V  A  $  �  �  l  W  7  �  �  �  �  �  �  �  `  D  C  G      �  �  �  �  �  �  �  �  T  F      A        
  	                                                             	return data          data['partnership']=partnership         partnership=frappe.db.sql("select MONTHNAME(creation) as Month, ifnull((select sum(amount) from `tabPartnership Record` where giving_or_pledge='Giving' and partnership_arms=p.partnership_arms and year(creation)=year(p.creation) and MONTH(creation)=MONTH(p.creation)),0) as `giving`,ifnull((select sum(amount) from `tabPartnership Record` where giving_or_pledge='Pledge' and partnership_arms=p.partnership_arms and year(creation)=year(p.creation) and MONTH(creation)=MONTH(p.creation)),0) as pledge,partnership_arms from `tabPartnership Record` p where creation between date_sub(now(),INTERVAL 120 day) and now() and  partnership_arms is not null group by year(creation), MONTH(creation),partnership_arms",as_dict=1)                  data['membership_strength']='0'         else:                data['membership_strength']=membership_strength         if membership_strength:         membership_strength=frappe.db.sql("select a.month,a.total_member_count,b.conversion as `new_converts` from ( SELECT COUNT(name) AS total_member_count,MONTHNAME(creation) as month FROM `tabMember` WHERE creation BETWEEN date_sub(now(),INTERVAL 90 day) AND now() GROUP BY YEAR(creation),MONTH(creation)) a, (select MONTHNAME(creation) as month ,count(ftv_id_no) as conversion from tabMember where ftv_id_no is not null group by YEAR(creation), MONTH(creation)) b where a.month=b.month",as_dict=1)          data['first_timers']=first_timers 	first_timers=frappe.db.sql("select a.`Week` as `Week3`,b.`Month` as `Month3`,c.`Year` as `Year3` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() ) a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b,(select count(name) as `Year` from `tabFirst Timer` where                      creation between date_sub(now(),INTERVAL 1 Year) and now())c" , as_dict=1)          data['new_converts']=new_born 	new_born=frappe.db.sql("select a.`Week` as `Week2`,b.`Month` as `Month2`,c.`Year` as `Year2` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() and is_new_born='Yes') a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now() and is_new_born='Yes') b,(select count(name)             as `Year` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Year) and now() and is_new_born='Yes')c" , as_dict=1)          data['invities_contacts']=new_visitor 	new_visitor=frappe.db.sql("select a.`Week` as `Week1`,b.`Month` as `Month1`,c.`Year` as `Year1` from (select count(name) as `Week` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 WEEK)  and now()) a,(select count(name) as `Month` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b, (select count(name) as `Year` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Year) and now())c", as_dict=1)          data['dates']=dates         dates['Year1']='Year : 2015'         dates['Month1']='Month : Sep'         dates['Week1']='Week : 2'  	dates={}         data={}             }                   "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def dashboard(data): @frappe.whitelist(allow_guest=True)        return ma.name+" created Successfully"     ma.insert(ignore_permissions=True)     ma = frappe.get_doc(dts)     del dts['name'] ad  !   �               �  �  �  �  �  �	  �	  �  �  S  D    >       �  �  Q  8    �  �    t  �   �   �   �                                             #data['invities_contacts']=new_visitor         #(select count(name) as `Year` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Year) and now())c", as_dict=1)         #and now()) a,(select count(name) as `Month` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b,\ 	#new_visitor=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 WEEK) \                 data['new_visitor']='0'         else:                 data['new_visitor']=new_visitor[0][0]         if new_visitor :         new_visitor=frappe.db.sql("select count(name) from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 WEEK) and now()")         # old code            #return data         #data['partnership']=partnership         #partnership=frappe.db.sql("select MONTHNAME(creation) as Month, ifnull((select sum(amount) from `tabPartnership Record` where giving_or_pledge='Giving' and partnership_arms=p.partnership_arms and year(creation)=year(p.creation) and MONTH(creation)=MONTH(p.creation)),0) as `giving`,ifnull((select sum(amount) from `tabPartnership Record` where giving_or_pledge='Pledge' and partnership_arms=p.partnership_arms and year(creation)=year(p.creation) and MONTH(creation)=MONTH(p.creation)),0) as pledge,partnership_arms from `tabPartnership Record` p where creation between date_sub(now(),INTERVAL 120 day) and now() and  partnership_arms is not null group by year(creation), MONTH(creation),partnership_arms",as_dict=1)         #        data['membership_strength']='0'         #else:         #        data['membership_strength']=membership_strength         #if membership_strength: 	#membership_strength=frappe.db.sql("select a.month,a.total_member_count,b.conversion as `new_converts` from ( SELECT COUNT(name) AS total_member_count,MONTHNAME(creation) as month FROM `tabMember` WHERE creation BETWEEN date_sub(now(),INTERVAL 90 day) AND now() GROUP BY YEAR(creation),MONTH(creation)) a, (select MONTHNAME(creation) as month ,count(ftv_id_no) as conversion from tabMember where ftv_id_no is not null group by YEAR(creation), MONTH(creation)) b where a.month=b.month",as_dict=1)         #data['first_timers']=first_timers         #first_timers=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() )         	a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b,(select count(name) as `Year` from `tabFirst Timer` where        		creation between date_sub(now(),INTERVAL 1 Year) and now())c" , as_dict=1) 	         #data['new_converts']=new_born         #new_born=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() and         	is_new_born='Yes') a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now() and is_new_born='Yes') b,(select count(name)         	as `Year` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Year) and now() and is_new_born='Yes')c" , as_dict=1)          #data['invities_contacts']=new_visitor         #new_visitor=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 WEEK)      and now()) a,(select count(name) as `Month` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b,      (select count(name) as `Year` from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 Year) and now())c", as_dict=1) ad     �      &       c  N      �  +  f  �  �  �      �  �  �  �
  
  �	  �	  �	  �  �  �  }  N  =  M  -  �  �  �  �  �  �  Q  C    �   �               	#partnership=frappe.db.sql("select MONTHNAME(creation) as Month, ifnull(sum(amount),0) as `giving`,ifnull(sum(amount),0) as pledge,partnership_arms from `tabPartnership Record` where creation between date_sub(now(),INTERVAL 120 day) and now() and  partnership_arms is not null group by year(creation), MONTH(creation),partnership_arm ",as_dict=1)                data['partnership']='0'         else:                data['partnership']=partnership         if partnership: 	partnership=frappe.db.sql("select MONTHNAME(creation) as Month, ifnull(sum(amount),0) as `giving`,ifnull(sum(amount),0) as pledge from `tabPartnership Record` where creation between date_sub(now(),INTERVAL 1 Year) and now() group by year(creation), MONTH(creation)",as_dict=1)         #partnership=frappe.db.sql("select MONTHNAME(creation) as Month, count(name) as `giving`,count(name) as pledge from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Year) and now() group by year(creation), MONTH(creation)",as_dict=1)                data['membership_strength']='0'         else:                data['membership_strength']=membership_strength         if membership_strength: 	membership_strength=frappe.db.sql("select a.month,a.total_member_count,b.conversion as `new_converts` from ( SELECT COUNT(name) AS total_member_count,MONTHNAME(creation) as month FROM `tabMember` WHERE creation BETWEEN date_sub(now(),INTERVAL 1 YEAR) AND now() GROUP BY YEAR(creation),MONTH(creation)) a, (select MONTHNAME(creation) as month ,count(ftv_id_no) as conversion from tabMember where ftv_id_no is not null group by YEAR(creation), MONTH(creation)) b where a.month=b.month",as_dict=1)         #membership_strength=frappe.db.sql("select MONTHNAME(creation) as Month, count(name) as `New Users`,count(name) as Revisited from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Year) and now() group by year(creation), MONTH(creation)",as_list=1)                data['visitor_last_months']='0'         else:                data['visitor_last_months']=visitor_last_months[0][0]         if visitor_last_months:         visitor_last_months=frappe.db.sql("select count(name) from `tabInvitees and Contacts` where creation between date_sub(now(),INTERVAL 1 WEEK) and now()")          #data['first_timers']=first_timers         #		creation between date_sub(now(),INTERVAL 1 Year) and now())c" , as_dict=1)         #	a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now()) b,(select count(name) as `Year` from `tabFirst Timer` where \ 	#first_timers=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() ) \                 data['first_timers']='0'         else:                 data['first_timers']=first_timers[0][0]         if first_timers:         first_timers=frappe.db.sql("select count(name) from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 YEAR) and now()") 	         #data['new_converts']=new_born         #	as `Year` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Year) and now() and is_new_born='Yes')c" , as_dict=1)         #	is_new_born='Yes') a,(select count(name) as `Month` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 Month) and now() and is_new_born='Yes') b,(select count(name) \ 	#new_born=frappe.db.sql("select a.`Week`,b.`Month`,c.`Year` from (select count(name) as `Week` from `tabFirst Timer` where creation between date_sub(now(),INTERVAL 1 WEEK) and now() and \                 data['new_born']='0'            else:                 data['new_born']=new_born[0][0]         if new_born:         new_born=frappe.db.sql("select count(name) from `tabMember` where creation between date_sub(now(),INTERVAL 1 YEAR) and now() and is_new_born='Yes'") ad  �  �     N       �  �  �  �  �  j  �  �  �  �  �  N  B  �  �  �  \  9     �  �  t  c  C    �  5  %  $  #  �
  �
  �
  G
  *
  
  
  �	  �	  �	  �  �  �  �  �  s  ]  >    �  i  H  2    �  �  �  �  ~  a  =    �  �  �  �  t  Y  7    �  �  �  �  �  y    �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    elif dts['search']=='Leader':                 qry="select church,pcf,senior_cell,name as cell from tabCells where "+cstr(key)+"='"+cstr(value)+"'"         if dts['search']=='Group':                 value=1                 key='1'         else:                 value=dts['region']                 key='region'         elif dts['region']:                 value=dts['zone']                 key='zone'         elif dts['zone']:                 key1='church_group'                 value=dts['group']                 key='group_church'         elif dts['group_church']:                 key1='church_name'                 value=dts['church']                 key='church'         if dts['church']:         qry=''             }                          "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data)         #frappe.response.update(frappe.sessions.get())         import frappe.sessions def search_glm(data): @frappe.whitelist(allow_guest=True)        return "The Partnership Record '" +cstr(dts['name'])+ "' Is updated successfully."     frappe.db.sql("update `tabPartnership Record` set giving_or_pledge='%s',amount='%s' where name='%s'" %(dts['giving_or_pledge'],dts['amount'],dts['name']) ,as_dict=True)         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def update_partnership_arm(data): @frappe.whitelist(allow_guest=True)       return data     data=frappe.db.sql("select name,partnership_arms,ministry_year,is_member,member,date,church,giving_or_pledge,amount from `tabPartnership Record`  where name='%s'" %(dts['name']) ,as_dict=True)         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def partnership_arm_details(data): @frappe.whitelist(allow_guest=True)      return data     data=frappe.db.sql("select name,church,partnership_arms,giving_or_pledge,sum(amount) as amount from `tabPartnership Record` group by church,giving_or_pledge ",as_dict=True)         }                   "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data) def partnership_arm(data): @frappe.whitelist(allow_guest=True)          return data         #data['partnership']=partnership ad     ^     K       9    w  p    �  �  �  �  �  z  ]  Q  :  �
  �
  �
  m
  M
  
   
  �	  Q	  �  �  �  j     �  �  t  G    �  �  �  �  �  �    �  �  �  �  i  [  9    �  �  �  �  �  �  j  R  5  �  �  }  h  H  	  �  �  �  �  �  h  K  �  �  �  ~  ^  ]                                        "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def list_members_details(data): @frappe.whitelist(allow_guest=True)  	return res         res=frappe.db.sql("select name from tabMember",as_dict=1)             }                 "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def list_members(data): @frappe.whitelist(allow_guest=True)               return ma.name             ma.insert(ignore_permissions=True)             ma = frappe.get_doc(rr)             del rr['password']             #del rr['name']         for rr in dts['records']:             }                 "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def member(data): @frappe.whitelist(allow_guest=True)          }             "comment": comment.as_dict()             "file_url": filedata.file_url,             "file_name": filedata.file_name,             "name": filedata.name,         return { 	#frappe.errprint(filedata.name,filedata.file_name,filedata.file_url,comment.as_dict())              frappe.db.sql("update tabMember set image=%s where name=%s",(filedata.file_url,dts['name'])) 	if dts['tbl']=='Member':              _("Added {0}").format("<a href='{file_url}' target='_blank'>{file_name}</a>".format(**filedata.as_dict())))         comment = frappe.get_doc(dts['tbl'], dts['name']).add_comment("Attachment",         filedata=save_file(fname=dts['filename'],content=base64.b64decode(dts['fdata']),dt=dts['tbl'],dn=dts['name'])         from frappe.utils.file_manager import  save_file             }                 "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	#frappe.errprint(dts) 	#print dts         dts=json.loads(data) def file_upload(data): @frappe.whitelist(allow_guest=True)          return data         data=frappe.db.sql(qry,as_dict=True)         #return qry 		 qry="select name , member_name, church,church_group,zone,region,phone_1,email_id from tabMember " 	else:                 qry="select name , member_name, church,church_group,zone,region,phone_1,email_id from tabMember where member_name like '%"+cstr(dts['member'])+"%'"         elif 'member' in dts:                 qry="SELECT ttl.church_name AS church,ttl.church_group AS group_type,ttl.member_name AS member_name,ttl.phone_no AS phone_no FROM ( SELECT cc.name AS church_name, cc.church_group AS church_group, mmbr.member_name AS member_name, mmbr.phone_1 AS phone_no, cc.zone As zone, cc.region as regin FROM tabChurches cc, ( SELECT m.member_name, m.phone_1, userrol.defvalue AS defvalue FROM tabMember m , ( SELECT a.name AS name, c.defvalue AS defvalue FROM tabUser a, tabUserRole b, tabDefaultValue c WHERE a.name=b.parent AND a.name=c.parent AND b.role='Church Pastor' AND c.defkey='Churches' ) userrol WHERE m.user_id=userrol.name) mmbr WHERE cc.name=mmbr.defvalue) ttl WHERE ttl."+key1+"='"+value+"'" ad  �   1     M       �  �  �  d  Y  F  E  !    �  i  H  2    �  �  �  9  #  �
  �
  �
  �
  �
  �
  
  �	  �	  �	  �	  \	  N	  $	  �  �  �  �  U  9  !  �  �  �  g  G  +    �  �  �  k  A    �  �  �  �  �  �  �  h  `  G  8    �  j  X  G  '  �  �  �    �  ;  1  0                                                                                                                                                                                                                                       else:        qry="select name,member_name as ftv_name,email_id,phone_1 from tabMember where email_id in (select u.name from tabUser u,tabUserRole ur where u.enabled=1 and ur.role='Member') "     elif dts['tbl']=='Member':        qry="select name,ftv_name ,email_id,phone_1 from `tabFirst Timer` where email_id in (select u.name from tabUser u,tabUserRole ur where u.enabled=1 and ur.role='Member' )"     if dts['tbl']=='FT':         }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     from frappe.model.db_query import DatabaseQuery     #print dts     dts=json.loads(data)     """     this will return recipents details     """ def message_braudcast_details(data): @frappe.whitelist(allow_guest=True)            return "Your profile updated successfully"         obj1.save(ignore_permissions=True)         obj1.new_password=dts['password'] 	obj1=frappe.get_doc('User',dts['username']) 	obj.save(ignore_permissions=True) 	obj.phone_1=dts['phone_1'] 	obj.experience_years=dts['experience_years'] 	obj.marital_info=dts['marital_info'] 	obj.phone_2=dts['phone_2'] 	obj.email_id2=dts['email_id2'] 	obj.member_name=dts['member_name'] 	obj.core_competeance=dts['core_competeance'] 	obj.educational_qualification=dts['educational_qualification'] 	obj.date_of_birth=dts['date_of_birth'] 	obj.image=dts['image'] 	obj.address=dts['address'] 	obj.employment_status=dts['employment_status'] 	obj.industry_segment=dts['industry_segment'] 	#obj.email_id=dts['email_id'] 	obj.office_address=dts['office_address'] 	obj.yearly_income=dts['yearly_income'] 	obj=frappe.get_doc('Member',dts['name'])             }                 "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def update_my_profile(data): @frappe.whitelist(allow_guest=True)          return res         res=frappe.db.sql(qr1,as_dict=1) 	#rappe.errprint(qr1)         qr1="select m.name,m.member_name,m.date_of_birth,m.phone_1,m.phone_2,m.email_id,m.email_id2,m.address,m.office_address,m.employment_status,m.industry_segment,m.yearly_income,m.experience_years,m.core_competeance,m.educational_qualification,null AS `password`,m.image,m.marital_info from tabMember m,tabUser u where m.email_id=u.name and u.name='"+dts['username']+"'"             }                 "message":"User name or Password is incorrect"                 "status":"401",             return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) def get_my_profile(data): @frappe.whitelist(allow_guest=True)          return res 	print res         res=frappe.db.sql(qr1,as_dict=1) 	qr1="select name,member_name,date_of_birth,phone_1,phone_2,email_id,email_id2,address,office_address,employment_status,industry_segment,yearly_income,experience_years,core_competeance,educational_qualification,null AS `password`,image,marital_info from tabMember where name='"+dts['name']+"'"             }                 "message":"User name or Password is incorrect" ad     �     l       �  �  �  �  �  _  Z  D  �  �  �  �  �  Q  M  F  <  �  �  
  �  P  .         �  �  �  �    s  U  I  �
  �
  �
  �
  z
  X
  
  
  �	  �	  �	  �	  n	  "	  !	   	  �  �  �  �  �  �  �    �  �  �  �  �  �  4    �  �  �  �  p  A    �  �  �  �  o  Z  +  �  �  �  �  �  �  b  J  E        �  �  w  ]  N  C  /  �  �  �  �  a      �  �  �                     		obj=frappe.new_doc("Cells") 	else:                 }                   "message":"You have no permission to create Senior Cell"                   "status":"403",                 return {         if not frappe.has_permission(doctype="Cells", ptype="create",user=dts['username']): 		} 		  "message":"User name or Password is incorrect" 		  "status":"401", 		return { 	if not valid: 	valid=frappe.db.sql(qry) 	qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	print data 	dts=json.loads(data) 	"""  	Need to check validation/ duplication  etc 	""" def create_cells(data): @frappe.whitelist(allow_guest=True)   		                 		return "Successfully created senior Cell '"+obj.name+"'" 		obj.insert(ignore_permissions=True) 		obj.contact_email_id=dts['contact_email_id'] 		obj.contact_phone_no=dts['contact_phone_no'] 		obj.pcf=dts['pcf'] 		obj.church=dts['church'] 		obj.church_group=dts['church_group'] 		obj.region=dts['region'] 		obj.zone=dts['zone'] 		obj.meeting_location=dts['meeting_location'] 		obj.senior_cell_code=dts['senior_cell_code'] 		obj.senior_cell_name=dts['senior_cell_name'] 		obj=frappe.new_doc("Senior Cells") 	else:                 }                   "message":"You have no permission to create Senior Cell"                   "status":"403",                 return {         if not frappe.has_permission(doctype="Senior Cells", ptype="create",user=dts['username']): 		} 		  "message":"User name or Password is incorrect" 		  "status":"401", 		return { 	if not valid: 	valid=frappe.db.sql(qry) 	qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	dts=json.loads(data) 	"""  	Need to check validation/ duplication  etc 	""" def create_senior_cells(data): @frappe.whitelist(allow_guest=True)                   return "Successfully updated device id '"+obj.device_id+"'" 		#print obj.device_id 		obj.save(ignore_permissions=True)                 obj.device_id=device_id 		obj=frappe.get_doc("User",username)         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry) 	#print qry         qry="select user from __Auth where user='"+cstr(username)+"' and password=password('"+cstr(userpass)+"') " 	#print dts         #dts=json.loads(data)         """          Need to check validation/ duplication  etc         """ def create_push_notification(device_id,username,userpass): @frappe.whitelist(allow_guest=True)   		return data 		data['user_values']=user_values 		#user_values=frappe.db.sql("select defkey,defvalue from `tabDefaultValue`  where parent=%(user)s", {"user":dts['username']},as_dict=True) 		user_values=frappe.db.sql(qry,as_dict=True) 		qry="select defkey,defvalue from `tabDefaultValue`  where defkey not like '_list_settings:%' and defkey not like '_desktop_items%' and parent='"+dts['username']+"'" 		data['roles']=roles 		roles=frappe.db.sql("select role from `tabUserRole` where parent=%(user)s", {"user":dts['username']},as_dict=True) 		data={} 	else: 		} 			"message":"User name or Password is incorrect" 			"status":"401", 		return { 	if not valid: 	valid=frappe.db.sql(qry) 	qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	dts=json.loads(data) 	""" 	Get user name and password from user and returns roles and its def key and defvalue 	""" def user_roles(data): @frappe.whitelist(allow_guest=True)  # gangadhar ad  7   �     c       �  �  �  r  M  6    �  �  �  �  f  @  8     �  �  �  �  �  �  �  �  q  e  H  �  �  �  w  U      �  �  k  '      �
  �
  �
  [
  0
  
  �	  �	  �	  :	  (	  	  	  �  �  �  �  �  h  �  �  �  �  u  4  "  �  �  �  G  5  '  �  �  �  p  E    �  �  �  Q  ?  $  #  �  �  �  {  H  C  &  �  �  n  U  3  �  �  �  �                                                                          }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) 	"""         Need to check validation/ duplication  etc 	No Need to send sms,push notification and email , it should be on attendence update on every user. 	""" def create_meetings(data): @frappe.whitelist(allow_guest=True)                  return ret                 }                         "message":"Successfully updated Event '"+obj.name+"'"                 ret={                 obj.save(ignore_permissions=True)                 obj.description=dts['description']                 obj.address=dts['address']                 obj.ends_on=dts['ends_on']                 obj.starts_on=dts['starts_on']                 obj.type=dts['type']                 obj.subject=dts['subject']                 obj=frappe.get_doc("Event",dts['name'])         else:                 }                   "message":"You have no permission to create Cell"                   "status":"403",                 return {         if not frappe.has_permission(doctype="Event", ptype="create",user=dts['username']):                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data)         """         Need to check validation/ duplication  etc         """ def update_event(data): @frappe.whitelist(allow_guest=True)                  return ret                 }                         "message":"Successfully created Event '"+obj.name+"'"                 ret={                 obj.insert(ignore_permissions=True)                 obj.description=dts['description']                 obj.address=dts['address']                 obj.ends_on=dts['ends_on']                 obj.starts_on=dts['starts_on']                 #obj.type=dts['type']                 obj.subject=dts['subject']                 obj=frappe.new_doc("Event")         else:                 }                   "message":"You have no permission to create Cell"                   "status":"403",                 return {         if not frappe.has_permission(doctype="Event", ptype="create",user=dts['username']):                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data)         """         Need to check validation/ duplication  etc         """ def create_event(data): @frappe.whitelist(allow_guest=True)    		return ret 		} 			"message":"Successfully created Cell '"+obj.name+"'" 		ret={ 		obj.insert(ignore_permissions=True) 		obj.contact_email_id=dts['contact_email_id'] 		obj.contact_phone_no=dts['contact_phone_no'] 		obj.pcf=dts['pcf'] 		obj.church=dts['church'] 		obj.church_group=dts['church_group'] 		obj.region=dts['region'] 		obj.zone=dts['zone'] 		obj.senior_cell=dts['senior_cell'] 		obj.address=dts['address'] 		obj.meeting_location=dts['meeting_location'] 		obj.cell_code=dts['cell_code'] 		obj.cell_name=dts['cell_name'] ad  b   �     \       �  �  x  -  !    �  �  �  �  �  �  �  �  '    �  �  �  y  1      �  �  �  g  >  7    �
  �
  �
  �
  Z
  =
  
  �	  �	  �	  �	  U	  G	  �  �  �  �  �  �  �  �  g  b  E  9  �  �  �  h  F    �  �  �  �  d  1    �  ~  J  6        �  �  �  �  �  �    �  �  �  �  T  B  4  �  �  �  �                                                                                                                    #data=frappe.db.sql("select name,member,member_name,present from `tabInvitation Member Details` where parent=%s",dts['meeting_id'],as_dict=True) 		#frappe.session.user=dts['username'] 		#frappe.local.session_obj = Session(user=dts['username'], resume=resume,full_name=dts['username'], user_type="System User")         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) 	""" 	Get all participents of selected meeting 	""" def meetings_members(data): @frappe.whitelist(allow_guest=True)                  return data 	       #print data                data=frappe.db.sql(qry,as_dict=True) 	       #print qry                qry="select name as meeting_name,meeting_subject , from_date as meeting_date ,venue from `tabAttendance Record` where 1=1 " 	       #print mcond 	       #mcond=get_match_cond("Attendance Record") 	       #print frappe.session.user 	       #print dts['username'] 	       from erpnext.controllers.queries import get_match_cond         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	#print dts         dts=json.loads(data) 	""" 	Need to add filter of permitted records for user 	""" def meetings_list(data): @frappe.whitelist(allow_guest=True)           return ret         }                         "message":"Successfully created Cell '"+obj.name+"'"         ret={ 	print "Successfully created Cell '"+obj.name+"'"         obj.insert(ignore_permissions=True)         obj.pcf=dts['pcf']         obj.church=dts['church']         obj.church_group=dts['church_group']         obj.region=dts['region']         obj.zone=dts['zone']         obj.senior_cell=dts['senior_cell']         obj.cell=dts['cell']         obj.venue=dts['venue']         obj.to_date=dts['to_date']         obj.from_date=dts['from_date'] 	        obj.meeting_sub=dts['meeting_sub'] 	else: 		obj.meeting_subject=dts['meeting_sub'] 	if dts['meeting_category']=="Cell Meeting":         obj.meeting_category=dts['meeting_category']         obj=frappe.new_doc("Attendance Record") 	#print data         #return "hello"                 }	                 "message":"To Date should be greater than From Date..!"                 "status":"402",                 return {             if dts['from_date'] >= dts['to_date']:         if dts['from_date'] and dts['to_date']:                 }                 "message":"Attendance Record is already created for same details on same date "                 "status":"401",             return {         if res:         res=frappe.db.sql("select name from `tabAttendance Record` where (cell='%s' or church='%s') and from_date like '%s%%' and to_date like '%s%%'"%(dts['cell'],dts['church'],f_date,t_date))         t_date=tdate[0]         tdate=dts['to_date'].split(" ")         f_date=fdate[0]         fdate=dts['from_date'].split(" ") 	#return "hello" 		        } 				"message":"You have no permission to create Meeting Attendance Record" 				"status":"403", 		        return { 	if not frappe.has_permission(doctype="Attendance Record", ptype="create",user=dts['username']): ad     S     K         �  �  �  �  �  �  S  N  1  %  �  �  m  T  2  �  �  �  �  U  �      �
  �
  �
  I
  	  	  �  r  F  E  D        �  �  �  �  ;      �  �  �  v  h  �  �  �  �  �  �  �  S  N  1  $  �  �  l  S  1  �  �  �  �  o  ;  �  x  w  S  R             @frappe.whitelist(allow_guest=True)                  return "Updated Attendance"                         frappe.db.sql("update `tabInvitation Member Details` set present=%s where name=%s",(record['present'],record['name']),debug=1)                                 record['present']=0                         if not record['present'] :                 for record in dts['records']:         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	#print(dts)         dts=json.loads(data) 	""" 	Member can mark their attandence of meeting 	""" def mark_my_attendance(data): @frappe.whitelist(allow_guest=True)                   return data                 data=frappe.db.sql("select a.name as meeting_name,a.meeting_category as meeting_category, a.meeting_subject as meeting_subject,a.from_date as from_date,a.to_date as to_date,a.venue as venue,b.name as name,ifnull(b.present,0) as present from `tabAttendance Record`  a,`tabInvitation Member Details` b where a.name=b.parent and b.email_id=%s",dts['username'],as_dict=True)         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "         dts=json.loads(data) 	""" 	Meeting list of member user 	""" def meetings_list_member(data): @frappe.whitelist(allow_guest=True)                   return "Updated Attendance" 				#	res = gcm.json_request(registration_ids=res[0], data=data,collapse_key='uptoyou', delay_while_idle=True, time_to_live=3600) 				#	print res[0] 				#	print reg_ids 				#	reg_ids=['APA91bGKibKhhg2RssK2eng8jXW7Gzhmq5_nDcxr8OiAxPSB62xlMdJdSPKCGO9mPF7uoLpT_8b-V0MdY33lc7fTNdh6U965YTQD3sIic_-sY3C45fF5dUEwVuVo8e2lmDduN4EUsHBH','APA91bHXuIe7c8JflytJnTdCOXlWzfJCM2yt5hGgwaqzIbNfGjANhqzLgrVCoSno70hKtygzg_W7WbE4lHeZD_LeQ6CSc_5AteGY1Gh6R7NXihVnE45K91DOPxgtnF5ncN4gSJYiX0_N'] 				#	data = {'param1': 'new attendance updated sussessfully ....'} 				#	gcm = GCM('AIzaSyBIc4LYCnUU9wFV_pBoFHHzLoGm_xHl-5k') 				#	from gcm import GCM 				#if res and dts['push']=='1': 				#print res 				res=frappe.db.sql("select device_id from tabUser where name=(select email_id from `tabInvitation Member Details` where name=%s) ",record['name'],as_list=True,debug=1)                                 frappe.db.sql("update `tabInvitation Member Details` set present=%s where name=%s",(record['present'],record['name']))                         if record['present']=='0' or record['present']=='1' :                 for record in dts['records']:         else:                 }                   "message":"User name or Password is incorrect"                   "status":"401",                 return {         if not valid:         valid=frappe.db.sql(qry)         qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	#print dts         dts=json.loads(data) 	""" 	Need to add provision to send sms,push notification and emails on present and absent 	""" def meetings_attendance(data): @frappe.whitelist(allow_guest=True)                   return data 		data=frappe.db.sql("select b.name,b.member,b.member_name,b.present,a.venue,a.meeting_subject,a.from_date from `tabAttendance Record` a,`tabInvitation Member Details` b  where a.name=b.parent and  a.name=%s",dts['meeting_id'],as_dict=True) ad     [     L       �  �  g  �  �  �  �  C  8  �  �  �  �  �  �  �  �  �  �  v  q  [  *  �  �  �  |  h  5  1  �
  
  �	  �	  �	  �	  �	  �  �  �  [    g  �  �  �  �  �  1  %  �  �  {  �  �  �  j  S    V  N  B    �  �  L  "  �  �  �  �  �  �  �    [  Z                 @frappe.whitelist(allow_guest=True)   	#	} 	#			"message":"No Records Found" 	#			"status":"200", 	#	return { 	#else: 	#	return frappe.db.sql("""select name from `tab%s` """%(dts['tbl']), as_dict=1) 	#elif ("System Manager" in user_roles ): 	#	return frappe.db.sql("""select name from `tab%s` where %s"""%(dts['tbl'], ' or '.join(match_conditions)), as_dict=1) 	#	cond = 'where ' + ' or '.join(match_conditions) 	#if match_conditions   : 	#user_roles = frappe.get_roles(dts['username']) 	#cond = '' 	##		)) 	##				or `tab{doctype}`.`{fieldname}` in ({values}))""".format(doctype=dts['tbl'],fieldname=df.fieldname,values=", ".join([('"'+v+'"') for v in user_permissions[df.options]]) 	##		match_conditions.append("""(ifnull(`tab{doctype}`.`{fieldname}`, "")="" 	##		#print df.options 	##	for df in meta.get_fields_to_check_permissions(doctypes): 	##	#print doctypes 	##for doctypes in user_permissions: 	#		match_conditions.append(""" {fieldname} is null or {fieldname} ='{values}'""".format(doctype=dts['tbl'],fieldname=res[0][0],values=item['defvalue']))         #	if res:	         #	res=frappe.db.sql(qry) 	#	qry="select fieldname from tabDocField where options='"+cstr(item['defkey'])+"' and parent='"+cstr(dts['tbl'])+"'" 	#    else: 	#    	match_conditions.append(""" name ='{values}'""".format(values=item['defvalue'])) 	#    if item['defkey']==dts['tbl']: 	#for item in user_permissions: 	 	#match_conditions = [] 	##user_permissions=frappe.db.sql("select defkey,defvalue from tabDefaultValue where parent=%s " ,dts['username'],as_dict=1)   	##user_permissions1 =frappe.db.sql("""select defkey,defvalue from tabDefaultValue where parent=%s and parenttype='User Permission'""", (dts['username']),as_dict=True) 	##user_permissions = frappe.defaults.get_user_permissions(dts['username']) 	#role_permissions = frappe.permissions.get_role_permissions(meta, dts['username']) 	#meta = frappe.get_meta(dts['tbl'])  	return frappe.db.sql("""select name ,%s as record_name  from `tab%s` where %s"""%(','.join([x[0] for x in colmns ]),dts['tbl'], ' or '.join(match_conditions)), as_dict=1) 	#return ','.join([x[0] for x in colmns ]) 	        cond =' 1=1'	 	else: 		cond =  ' or '.join(match_conditions)      	if match_conditions   :     	colmns=frappe.db.sql("select fieldname from tabDocField where fieldtype !='Section Break' and fieldtype !='Column Break' and parent='%s' and fieldname like '%%_name%%' order by idx limit 6 " %(dts['tbl']),as_list=1 ) 	match_conditions=get_match_conditions(dts['tbl'],dts['username']) 		} 				"message":"User name or Password is incorrect" 				"status":"401", 		return { 	if not valid: 	valid=frappe.db.sql(qry) 	qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') " 	from frappe.model.db_query import DatabaseQuery 	dts=json.loads(data) 	""" 	Member can mark their attandence of meeting 	""" def get_masters(data): @frappe.whitelist(allow_guest=True)   	return match_conditions 			match_conditions.append(""" {fieldname} is null or {fieldname} ='{values}'""".format(doctype=doctype,fieldname=res[0][0],values=item['defvalue']))         	if res:	         	res=frappe.db.sql(qry) 		qry="select fieldname from tabDocField where options='"+cstr(item['defkey'])+"' and parent='"+cstr(doctype)+"'" 	    else: 	    	match_conditions.append(""" name ='{values}'""".format(values=item['defvalue'])) 	    if item['defkey']==doctype: 	for item in user_permissions: 	match_conditions = []	 	user_permissions=frappe.db.sql("select defkey,defvalue from tabDefaultValue where parent=%s ",username,as_dict=1)   	role_permissions = frappe.permissions.get_role_permissions(meta, username) 	meta = frappe.get_meta(doctype) def get_match_conditions(doctype,username): ad     �     Z       �  �  �  �  �  u  �  �  �  �  �  Y  K  �  h  X  /        �  �  �  �  �  �  	  �  �  �  �  j  Y  k
  [
  J
  I
  %
  	
  
  �	  �	  �	  �	  	  	  �  �  �  �  c  Y  Q  0       �  �  B  �  �  �  �  p  `  J    �  S  3  2    �  �  �  �  �  9    
  �  �  �  �  �  �  �  �  �  �  �                       def my_event_attendance(data): @frappe.whitelist(allow_guest=True)      return data                          where a.name=b.event_name and b.name=c.parent and c.id in (select a.name from tabMember a,tabUser b where a.email_id=b.name and b.name=%s) ",dts['username'],as_dict=True)     data=frappe.db.sql("select a.subject ,a.starts_on as event_date, a.address,c.name,c.person_name,ifnull(c.present,0) as present,comments from `tabEvent` a, `tabEvent Attendance` b,`tabEvent Attendace Details` c \         }                        "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data)     """     Member Event list     """ def my_event_list(data): @frappe.whitelist(allow_guest=True)      return "Updated Attendance" 		res = gcm.json_request(registration_ids=res[0], data=data,collapse_key='uptoyou', delay_while_idle=True, time_to_live=3600) 		data = {'param1': 'event attendance updated sussessfully ....'} 		gcm = GCM('AIzaSyBIc4LYCnUU9wFV_pBoFHHzLoGm_xHl-5k') 		from gcm import GCM 		#print res[0] 	if res and dts['push']=='1': 	#print res 	res=frappe.db.sql(qry,as_list=True) 	#print qry 	qry="select device_id from tabUser where name=(select email_id from tabMember where name='"+cstr(record['name'])+"')"         frappe.db.sql("update `tabEvent Attendace Details` set present=%s where id=%s",(record['present'],record['name']))             record['present']=0         if not record['present'] : 	#return record 	#frappe.errprint(type(record))     for record in dts['record']:                 }                 "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     #print dts     dts=json.loads(data)     """     update Event attendance     Give provisin for sms email and push notification     """ def event_attendance(data): @frappe.whitelist(allow_guest=True)                       return data     data=frappe.db.sql("select a.id as `name` ,a.person_name,ifnull(a.present,0) as present,a.comments from `tabEvent Attendace Details`  a,`tabEvent Attendance` b  where a.parent=b.name and b.event_name=%s",dts['event_id'],as_dict=True)         }                        "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     dts=json.loads(data)     """     Event details og selected event     """ def event_participents(data): @frappe.whitelist(allow_guest=True)               return data     data=frappe.db.sql(qry,as_dict=True)     #return qry     qry=" select name as event_name,address,starts_on as event_date,subject from tabEvent where "+get_permission_query_conditions(dts['username'])     from frappe.desk.doctype.event.event import get_permission_query_conditions         }                     "message":"User name or Password is incorrect"                 "status":"401",         return {     if not valid:     valid=frappe.db.sql(qry)     qry="select user from __Auth where user='"+cstr(dts['username'])+"' and password=password('"+cstr(dts['userpass'])+"') "     from frappe.model.db_query import DatabaseQuery     dts=json.loads(data)     """     Event List for user     """ def event_list(data): 